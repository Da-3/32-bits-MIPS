library ieee ; 
use ieee.std_logic_1164.all ;

entity top_level_entity is 
port ( 
		
		clk		: in 	std_logic;
		start		: in	std_logic;
		hit		: out std_logic
		

		
		);
		
end top_level_entity ; 

 architecture behav of top_level_entity is 
 begin 
 
 
 
 end behav;