library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CACHE_RAM is
	port(
		pc,data_in: 	in 	std_logic_vector(31 downto 0);
		ce,re,we:		in		std_logic;	
		data_out:		out	std_logic_vector(31 downto 0)
	);
end entity;


architecture rtl of CACHE_RAM is

type mem_array is array(0 to 127) of 
        std_logic_vector(31 downto 0);

signal mem: mem_array:=(
--R type without dependencies:
		--"00000001101101010100000000100000",  --add $t0,$t5,$s5
		--"00000001101101010100000000100010",  --sub $t0,$t5,$s5
		--"00000001101101010100000000100100",  --and $t0,$t5,$s5

--R type with RF dependency:
		--"00000001101101010100000000100000",    -- add $t0,$t5,$s5
		--"00000001101101010100100000100010",    -- sub $t1,$t5,$s5
		--"00000001101101010101000000100000",    -- add $t2,$t5,$s5
		--"00000001000101010101100000100100",    -- and $t3,$t0,$s5
		--"00000001000101010100000000100000",    -- add $t0,$t0,$s5

--R type with RAW dependencies: forwarding from MEM and WB to EXE stage

		--"00000001101101010100000000100000",    -- add $t0,$t5,$s5
		--"00000001000101010100100000100010",    -- sub $t1,$t0,$s5
		--"00000001101010000101000000100000",    -- add $t2,$t5,$t0
		--"00000001000101010101100000100100",    -- and $t3,$t0,$s5

--I,J type instructions without dependencies
		
		"10001100101010000000000000000000",     -- LW $t0, 0($R5)
		"00000000000000000000000000000000",     -- NOP
		"00100001000010000000000000000001",     -- addi $t0,$t0,1
		"10101100101010000000000000000000",     -- SW $t0, 0($R5)
		"00100000101001011111111111111111",     -- addi $R5,$R5,-1
		"00010000000001010000000000000010",     -- beq $zero, $R5, +2
		"00001000000000000000000000000000",     -- jump 0


		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000"
  );
--signal temp : std_logic_vector(31 downto 0);


begin

-- ce : input_enable (chip select)
-- re : read_enable
-- we	: write_enable

process(pc,data_in,ce,re,we) 
    begin
		if (ce = '1' and we = '1') then
			 mem(to_integer(unsigned(pc))) <= data_in;
		end if;
    end process;
	data_out <= mem(to_integer(unsigned(pc)));
end rtl;


